module ALU(
			input [2:0]					A,B,
			input [1:0]					Sel,
			output[4:0]					Out,
			output reg [4:0] 			result,
			output reg [13:0]			z
			);

	wire[4:0] temp;
	assign Out = result;
	
	always
	begin
		case (Sel)
		2'b00: result = A+B;
		2'b01: result = A-B;
		2'b10: result = A^B;
		2'b11: result = A<<1;
		
		endcase
		
		
		
		case (result[4:0])
		
		5'b00000 :
		z = 14'b10000001000000;					//Hex 0
		
		5'b00001 :
		z = 14'b10000001111001;					//Hex 1
		
		5'b00010 :
		z = 14'b10000000100100;					//Hex 2
		
		5'b00011 :
		z = 14'b10000000110000;					//Hex 3
		
		5'b00100 :
		z = 14'b10000000011001;					//Hex 4
		
		5'b00101 :
		z = 14'b10000000010010;					//Hex 5
		
		5'b00110 :
		z = 14'b10000000000010;					//Hex 6
		
		5'b00111 :
		z = 14'b10000001111000;					//Hex 7
		
		5'b01000 :
		z = 14'b10000000000000;					//Hex 8
		
		5'b01001 :
		z = 14'b10000010010000;					//Hex 9
		
		5'b01010 :
		z = 14'b11110011000000;					//Hex 10
		
		5'b01011 :
		z = 14'b11110011111001;					//Hex 11
		
		5'b01100 :
		z = 14'b11110010100100;					//Hex 12
		
		5'b01101 :
		z = 14'b11110010110000;					//Hex 13
		
		5'b01110 :
		z = 14'b11110010011001;					//Hex 14
		
		5'b01111 :
		z = 14'b11110010010010;					//Hex 15
		
		//subtraction
		
		5'b11111 :
		z = 14'b01111111111001;					//dec -1
				
		5'b11110 :
		z = 14'b01111110100100;					//dec -2
				
		5'b11101 :
		z = 14'b01111110110000;					//dec -3
				
		5'b11100 :
		z = 14'b01111110011001;					//dec -4
				
		5'b11011 :
		z = 14'b01111110010010;					//dec -5
				
		5'b11010 :
		z = 14'b01111110000010;					//dec -6
				
		5'b11001:
		z = 14'b01111111111000;					//dec -7
				
		5'b11000 :
		z = 14'b01111110000000;					//dec -8
		
		endcase
		
	end
	
endmodule
		
		
		
		
		


